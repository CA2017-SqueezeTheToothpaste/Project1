module Eq
(
	
);